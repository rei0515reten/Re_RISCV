module alu(input logic [31:0] SrcA,
	input logic [31:0] SrcB,
	input logic [2:0] ALUControl,
	input logic Zero,
	output logic [31:0] ALUResult);

	

endmodule
